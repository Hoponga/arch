////
//// Internal signal constants
////

// ALU
`define ALU_ADD      4'b0000
`define ALU_ADDU     4'b0001
`define ALU_SUB      4'b0010
`define ALU_SUBU     4'b0011 
`define ALU_AND      4'b0100 
`define ALU_OR       4'b0101  
`define ALU_XOR      4'b0110
`define ALU_NOR      4'b0111
`define ALU_SLT      4'b1000


`define R_TYPE       2'b00
`define I_TYPE       2'b01 
`define J_TYPE       2'b10



