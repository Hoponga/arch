/*
 *
 * Redistributions of any form whatsoever must retain and/or include the
 * following acknowledgment, notices and disclaimer:
 *
 * This product includes software developed by Carnegie Mellon University. 
 *
 * Copyright (c) 2004 by Babak Falsafi and James Hoe,
 * Computer Architecture Lab at Carnegie Mellon (CALCM), 
 * Carnegie Mellon University.
 *
 * This source file was written and maintained by Jared Smolens 
 * as part of the Two-Way In-Order Superscalar project for Carnegie Mellon's 
 * Introduction to Computer Architecture course, 18-447. The source file
 * is in part derived from code originally written by Herman Schmit and 
 * Diana Marculescu.
 *
 * You may not use the name "Carnegie Mellon University" or derivations 
 * thereof to endorse or promote products derived from this software.
 *
 * If you modify the software you must place a notice on or within any 
 * modified version provided or made available to any third party stating 
 * that you have modified the software.  The notice shall include at least 
 * your name, address, phone number, email address and the date and purpose 
 * of the modification.
 *
 * THE SOFTWARE IS PROVIDED "AS-IS" WITHOUT ANY WARRANTY OF ANY KIND, EITHER 
 * EXPRESS, IMPLIED OR STATUTORY, INCLUDING BUT NOT LIMITED TO ANYWARRANTY 
 * THAT THE SOFTWARE WILL CONFORM TO SPECIFICATIONS OR BE ERROR-FREE AND ANY 
 * IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE, 
 * TITLE, OR NON-INFRINGEMENT.  IN NO EVENT SHALL CARNEGIE MELLON UNIVERSITY 
 * BE LIABLE FOR ANY DAMAGES, INCLUDING BUT NOT LIMITED TO DIRECT, INDIRECT, 
 * SPECIAL OR CONSEQUENTIAL DAMAGES, ARISING OUT OF, RESULTING FROM, OR IN 
 * ANY WAY CONNECTED WITH THIS SOFTWARE (WHETHER OR NOT BASED UPON WARRANTY, 
 * CONTRACT, TORT OR OTHERWISE).
 *
 */

//////
////// MIPS 447: A single-cycle MIPS ISA simulator
//////

// Include the MIPS constants
`include "mips_defines.vh"
`include "internal_defines.vh"

////
//// The MIPS standalone processor module
////
////   clk          (input)  - The clock
////   inst_addr    (output) - Address of instruction to load
////   inst         (input)  - Instruction from memory
////   inst_excpt   (input)  - inst_addr not valid
////   mem_addr     (output) - Address of data to load
////   mem_data_in  (output) - Data for memory store
////   mem_data_out (input)  - Data from memory load
////   mem_write_en (output) - Memory write mask
////   mem_excpt    (input)  - mem_addr not valid
////   halted       (output) - Processor halted
////   reset        (input)  - Reset the processor
////   

module mips_core(/*AUTOARG*/
   // Outputs
   inst_addr, mem_addr, mem_data_in, mem_write_en, halted,
   // Inputs
   clk, inst_excpt, mem_excpt, inst, mem_data_out, rst_b
   );
   
   parameter text_start  = 32'h00400000; /* Initial value of $pc */

   // Core Interface
   input         clk, inst_excpt, mem_excpt;
   output [29:0] inst_addr;
   output [29:0] mem_addr;
   input  [31:0] inst, mem_data_out;
   output [31:0] mem_data_in;
   output [3:0]  mem_write_en;
   output        halted;
   input         rst_b;

   // Forced interface signals -- required for synthesis to work OK.
   // This is probably not what you want!
   

   // Internal signals
   wire [31:0] nextpc, branch_pc; 
   wire [31:0]   pc, nextnextpc, jump_target, branchtarget;
   wire [2:0] pc_src; 
   wire          exception_halt, syscall_halt, internal_halt;
   wire          load_epc, load_bva, load_bva_sel;
   wire [31:0]   rt_data, rs_data, rd_data, alu__out, r_v0;
   wire [31:0]   epc, cause, bad_v_addr;
   wire [4:0]    cause_code;
   wire [3:0]    alu_flags; 

   // Decode signals
   wire [31:0]   dcd_se_imm, dcd_se_offset, dcd_e_imm, dcd_se_mem_offset;
   wire [5:0]    dcd_op, dcd_funct2;
   wire [4:0]    dcd_rs, dcd_funct1, dcd_rt, dcd_rd, dcd_shamt;
   wire [15:0]   dcd_offset, dcd_imm;
   wire [25:0]   dcd_target;
   wire [19:0]   dcd_code;
   wire          dcd_bczft, imm_sign, is_shift;
   wire [1:0]    ins_type; 
   wire [4:0]    regfile_write_addr; 
   wire [31:0]   regfile_write_data; 
   wire [31:0]   alu_input_2; 
   wire [31:0]   imm_extend; 
   wire [31:0]   alu_input_1; 
   wire [2:0]    mem_read_bytes, mem_write_bytes; // how many bytes to read from/write to memory -- don't care if not a load/store instruction 
   
   // PC Management
   register #(32, text_start) PCReg(pc, nextpc, clk, ~internal_halt, rst_b);
   // register #(32, text_start+4) PCReg2(nextpc, nextnextpc, clk,
   //                                     ~internal_halt, rst_b);
   assign        inst_addr = pc[31:2];

   // Instruction decoding
   assign        dcd_op = inst[31:26];    // Opcode
   assign        dcd_rs = inst[25:21];    // rs field
   assign        dcd_rt = inst[20:16];    // rt field
   assign        dcd_rd = inst[15:11];    // rd field
   assign        dcd_shamt = inst[10:6];  // Shift amount
   assign        dcd_bczft = inst[16];    // bczt or bczf?
   assign        dcd_funct1 = inst[4:0];  // Coprocessor 0 function field
   assign        dcd_funct2 = inst[5:0];  // funct field; secondary opcode
   assign        dcd_offset = inst[15:0]; // offset field
        // Sign-extended offset for branches
   assign        dcd_se_offset = { {14{dcd_offset[15]}}, dcd_offset, 2'b00 };
        // Sign-extended offset for load/store
   assign        dcd_se_mem_offset = { {16{dcd_offset[15]}}, dcd_offset };
   assign        dcd_imm = inst[15:0];        // immediate field
   assign        dcd_e_imm = { 16'h0, dcd_imm };  // zero-extended immediate
        // Sign-extended immediate
   assign        dcd_se_imm = { {16{dcd_imm[15]}}, dcd_imm };
   assign        dcd_target = inst[25:0];     // target field
   assign        dcd_code = inst[25:6];       // Breakpoint code

   // synthesis translate_off
   always @(posedge clk) begin
     // useful for debugging, you will want to comment this out for long programs
     if (rst_b) begin
       $display ( "=== Simulation Cycle %d ===", $time );
       $display ( "[pc=%x, inst=%x] [op=%x, rs=%d, rt=%d, rd=%d, imm=%x, f2=%x] [reset=%d, halted=%d]",
                   pc, inst, dcd_op, dcd_rs, dcd_rt, dcd_rd, dcd_imm, dcd_funct2, ~rst_b, halted);
       $display ("[ctrl_we=%d, rd_data = %d, alu_out = %x, alu_flags = %b, imm_extend = %d, rt_data = %d]", ctrl_we, rd_data, alu__out, alu_flags, imm_extend, 
                   rt_data, mem_to_reg); 
       $display ("[mem_to_reg = %d, mem_addr = %x, mem_data_in = %x, mem_data_out = %x, regfile_write_data = %x, mem_excpt = %d]", 
                  mem_to_reg, mem_addr, mem_data_in, mem_data_out, regfile_write_data, mem_excpt); 
       $display ("[branch_result = %d, nextpc = %x, nextnextpc = %x, pc_src = %d, jumptarget = %x, branchtarget = %x]", 
                  branch_result, nextpc, nextnextpc, pc_src, jump_target, branchtarget);
     end
   end
   // synthesis translate_on

   // Let Verilog-Mode pipe wires through for us.  This is another example
   // of Verilog-Mode's power -- undeclared nets get AUTOWIREd up when we
   // run 'make auto'.
   
   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire [3:0]		alu__sel;		// From Decoder of mips_decode.v
   wire			ctrl_RI;		// From Decoder of mips_decode.v
   wire			ctrl_Sys;		// From Decoder of mips_decode.v
   wire			ctrl_we;		// From Decoder of mips_decode.v
   wire mem_to_reg;     // From Decoder of mips_decode.v 
   
   // End of automatics

   // Generate control signals
   mips_decode Decoder(/*AUTOINST*/
		       // Outputs
		       .ctrl_we		(ctrl_we),
		       .ctrl_Sys	(ctrl_Sys),
		       .ctrl_RI		(ctrl_RI),
		       .alu__sel	(alu__sel[3:0]),
           .alu__src  (alu__src), 
           .mem_to_reg(mem_to_reg),
           .ins_type(ins_type),
           .imm_sign(imm_sign),
           .is_shift(is_shift),
           .mem_read_bytes(mem_read_bytes),
           .mem_write_en(mem_write_en), 
           .mem_write_bytes(mem_write_bytes),

		       // Inputs
		       .dcd_op		(dcd_op[5:0]),
		       .dcd_funct2	(dcd_funct2[5:0]));
 
   // Register File
   // Instantiate the register file from reg_file.v here.
   // Don't forget to hookup the "halted" signal to trigger the register dump 
   assign regfile_write_addr = (ins_type == `J_TYPE && ctrl_we) ? 'hffffffff : (ins_type == `I_TYPE) ? dcd_rt : dcd_rd; 
   assign regfile_write_data = (ins_type == `J_TYPE && ctrl_we) ? (pc + 4) : (mem_to_reg) ? mem_data_out : alu__out; 

   

   regfile RegisterFile(
    .rs_num(dcd_rs), 
    .rt_num(dcd_rt), 
    .rd_num(regfile_write_addr), 
    .rd_data(regfile_write_data), 
    .rd_we(ctrl_we), 
    .clk(clk), 
    .rst_b(rst_b),
    .halted(halted), 
    .rs_data(rs_data), 
    .rt_data(rt_data)

   ); 

   // Execute
   assign imm_extend = (is_shift) ? dcd_shamt : (imm_sign) ? dcd_se_imm : dcd_e_imm; 

   assign alu_input_1 = (is_shift) ? dcd_shamt : rs_data; 

   assign alu_input_2 =(mem_to_reg) ? dcd_se_mem_offset : (alu__src) ? imm_extend : rt_data; 
   mips_ALU ALU(.alu__out(alu__out), 
                .alu__op1(alu_input_1),
                .alu__op2(alu_input_2),
                .alu__sel(alu__sel),
                .alu_flags(alu_flags));

   assign branch_result = ((dcd_op == `OP_BEQ) && alu_flags[3] == 1) || ((dcd_op == `OP_BNE) && alu_flags[3] != 1); 
   

   assign        mem_addr = (mem_to_reg) ? (alu__out[29:0] >> 2) : 0;
   assign        mem_data_in = rt_data;



   assign jump_target = {pc[31:28], dcd_target, 2'b00}; 
   assign branchtarget = pc + 4 + dcd_se_offset; 
   // assign nextnextpc = nextpc + 4; 
   assign branch_pc = (branch_result) ? branchtarget : pc + 4; 



   assign nextpc = (pc_src == 3'b1) ? jump_target : 
                   (pc_src == 3'b11 && branch_result == 1'b1) ? branchtarget : 
                        pc + 4;
   assign nextnextpc = (pc_src == 3'b1) ? jump_target + 4 : 
                   (pc_src == 3'b11 && branch_result == 1'b1) ? branchtarget + 4: 
                        nextpc + 4; 

   assign pc_src = (ins_type == `J_TYPE) ? 3'b1 : (ins_type == `B_TYPE) ? 3'b11 : 3'b0; 


   // // this block is basically our pc_sel mux 
   // always @(*) begin 
   //    case (pc_src) 
   //       3'b1: // jump instruction 
   //          nextpc = jump_target; 
   //       3'b11:   // branch instruction 
   //          nextpc = (branch_result) ? branchtarget : nextpc; 
   //    endcase 
      
   // end


 

   
   // Miscellaneous stuff (Exceptions, syscalls, and halt)
   exception_unit EU(.exception_halt(exception_halt), .pc(pc), .rst_b(rst_b),
                     .clk(clk), .load_ex_regs(load_ex_regs),
                     .load_bva(load_bva), .load_bva_sel(load_bva_sel),
                     .cause(cause_code),
                     .IBE(inst_excpt),
                     .DBE(1'b0),
                     .RI(ctrl_RI),
                     .Ov(1'b0),
                     .BP(1'b0),
                     .AdEL_inst(pc[1:0]?1'b1:1'b0),
                     .AdEL_data(1'b0),
                     .AdES(1'b0),
                     .CpU(1'b0));

   assign r_v0 = 32'h0a; // Good enough for now. To support syscall for real,
                         // you should read the syscall
                         // argument from $v0 of the register file 

   syscall_unit SU(.syscall_halt(syscall_halt), .pc(pc), .clk(clk), .Sys(ctrl_Sys),
                   .r_v0(r_v0), .rst_b(rst_b));
   assign        internal_halt = exception_halt | syscall_halt;
   register #(1, 0) Halt(halted, internal_halt, clk, 1'b1, rst_b);
   register #(32, 0) EPCReg(epc, pc, clk, load_ex_regs, rst_b);
   register #(32, 0) CauseReg(cause,
                              {25'b0, cause_code, 2'b0}, 
                              clk, load_ex_regs, rst_b);
   register #(32, 0) BadVAddrReg(bad_v_addr, pc, clk, load_bva, rst_b);

endmodule // mips_core


////
//// mips_ALU: Performs all arithmetic and logical operations
////
//// out (output) - Final result
//// in1 (input)  - Operand modified by the operation
//// in2 (input)  - Operand used (in arithmetic ops) to modify in1
//// sel (input)  - Selects which operation is to be performed

module mips_ALU(alu__out, alu_flags, alu__op1, alu__op2, alu__sel);

   output reg [31:0] alu__out;
   output reg [3:0] alu_flags; // from MSB to LSB, is Z C N V 
   input [31:0]  alu__op1, alu__op2;
   input [3:0]   alu__sel;
   wire set_ovflow; 
   wire pre_sign; 
   wire keep_sign_on_ovflow; 
   reg carry, zero; 

   assign pre_sign = alu__op1[31]; 
   
   
   // weird flag creation for N -- https://zipcpu.com/zipcpu/2017/08/11/simple-alu.html 
   assign keep_sign_on_ovflow = ((alu__sel == `ALU_ADD) && (alu__op1[31] == alu__op2[31])) || ((alu__sel == `ALU_SUB && (alu__op1[31] != alu__op2[31]))); 
   always @(*) begin 
      zero = ~|{alu__out  ^ 32'h00000000};
      $display("%b %b %d %d", alu__out, zero, alu__op1, alu__op2);
      alu_flags = {zero, carry, alu__out[31] ^ ((keep_sign_on_ovflow) && (pre_sign != alu__out[31])), 1'b0};
   end 
   always @(*) begin 
      
      case (alu__sel)
         `ALU_ADD: 
            {carry, alu__out} = alu__op1 + alu__op2; 
         `ALU_ADDU: 
            alu__out = alu__op1 + alu__op2; // right now, don't care about distinctions between unsigned and signed 
         `ALU_SUB: 
            {carry, alu__out} = alu__op1 - alu__op2; 
         `ALU_SUBU: 
            alu__out = alu__op1 - alu__op2; 
         `ALU_AND: 
            alu__out = alu__op1 & alu__op2; 
         `ALU_OR: 
            alu__out = alu__op1 | alu__op2; 
         `ALU_XOR: 
            alu__out = alu__op1 ^ alu__op2; 
         `ALU_SRL: 
            alu__out = alu__op2 >> alu__op1; 
         `ALU_SRA: 
            alu__out = alu__op2 >>> alu__op1; 
         `ALU_SLL: 
            alu__out = alu__op2 << alu__op1; 
         default: 
            {carry, alu__out} = alu__op1 + alu__op2; 

      endcase 
   end 

endmodule


//// register: A register which may be reset to an arbirary value
////
//// q      (output) - Current value of register
//// d      (input)  - Next value of register
//// clk    (input)  - Clock (positive edge-sensitive)
//// enable (input)  - Load new value?
//// reset  (input)  - System reset
////
module register(q, d, clk, enable, rst_b);

   parameter
            width = 32,
            reset_value = 0;

   output [(width-1):0] q;
   reg [(width-1):0]    q;
   input [(width-1):0]  d;
   input                 clk, enable, rst_b;

   always @(posedge clk or negedge rst_b)
     if (~rst_b)
       q <= reset_value;
     else if (enable)
       q <= d;

endmodule // register


////
//// adder
////
//// out (output) - adder result
//// in1 (input)  - Operand1
//// in2 (input)  - Operand2
//// sub (input)  - Subtract?
////
module adder(out, in1, in2, sub);
   output [31:0] out;
   input [31:0]  in1, in2;
   input         sub;

   assign        out = sub?(in1 - in2):(in1 + in2);

endmodule // adder


////
//// add_const: An adder that adds a fixed constant value
////
//// out (output) - adder result
//// in  (input)  - Operand
////
module add_const(out, in);

   parameter add_value = 1;

   output   [31:0] out;
   input    [31:0] in;

   assign   out = in + add_value;

endmodule // adder

// Local Variables:
// verilog-library-directories:("." "../447rtl")
// End:
